library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_pingpong is
end tb_pingpong;

architecture Behavioral of tb_pingpong is
    component pingpong is
        port(
            i_clk            : in STD_LOGIC;
            i_rst            : in STD_LOGIC;
            i_left_button    : in STD_LOGIC; 
            i_right_button   : in STD_LOGIC;
            i_speed_switch   : in STD_LOGIC;
            o_count          : out STD_LOGIC_VECTOR(7 downto 0)     
        );   
    end component;
    
    signal i_clk            : STD_LOGIC := '0';
    signal i_rst            : STD_LOGIC := '1';
    signal i_left_button    : STD_LOGIC := '0';
    signal i_right_button   : STD_LOGIC := '0';
    signal i_speed_switch   : STD_LOGIC := '0';
    signal o_count          : STD_LOGIC_VECTOR(7 downto 0);
    
    constant clk_period     : time := 10 ns;
    signal test_done        : boolean := false;
    
begin
    uut: pingpong
        port map (
            i_clk          => i_clk,
            i_rst          => i_rst,
            i_left_button  => i_left_button,
            i_right_button => i_right_button,
            i_speed_switch => i_speed_switch,
            o_count        => o_count
        );
    
    -- �����ͦ�
    clk_process: process
    begin
        while not test_done loop
            i_clk <= '0';
            wait for clk_period/2;
            i_clk <= '1';
            wait for clk_period/2;
        end loop;
        wait;
    end process;
    
    -- ���ը�E
    stim_proc: process
    begin
        -- Reset
        i_rst <= '0';
        wait for 100 ns;
        i_rst <= '1';
        wait for 100 ns;
        
        -- Test 1: �k�o�y�A�����~�]�k�o���^
        report "Test 1: Right serves, Left misses";
        i_right_button <= '1';
        wait for 100 ns;
        i_right_button <= '0';
        wait for 2000 ns;  -- ���ݲy���ʡA���䥢�~
        
        -- Test 2: ���o�y�A�k���~�]���o���^
        report "Test 2: Left serves, Right misses";
        i_left_button <= '1';
        wait for 100 ns;
        i_left_button <= '0';
        wait for 2000 ns;
        
        -- Test 3: ����若 - �k�o�y�A�Ӧ^�X���ᥪ���~
        report "Test 3: Rally with multiple hits";
        
        -- �k��o�y
        report "Right serves";
        i_right_button <= '1';
        wait for 50 ns;
        i_right_button <= '0';
        
        -- ���ݲy���ʨ�̥���]10000000�^
        wait until o_count = "10000000";
        wait for 10 ns;  -- �p����T�Oí�w
        report "Ball reached left side";
        
        -- �������y
        i_left_button <= '1';
        wait for 50 ns;
        i_left_button <= '0';
        
        -- ���ݲy���ʨ�̥k��]00000001�^
        wait until o_count = "00000001";
        wait for 10 ns;
        report "Ball reached right side";
        
        -- �k�����y
        i_right_button <= '1';
        wait for 50 ns;
        i_right_button <= '0';
        
        -- ���ݲy���ʨ�̥���]10000000�^
        wait until o_count = "10000000";
        wait for 10 ns;
        report "Ball reached left side again";
        
        -- �������y
        i_left_button <= '1';
        wait for 50 ns;
        i_left_button <= '0';
        
        -- ���ݲy���ʨ�̥k��]00000001�^
        wait until o_count = "00000001";
        wait for 10 ns;
        report "Ball reached right side again";
        
        -- �k�䤣���y�A���~
        report "Right misses - Left scores!";
        wait for 2000 ns;
        
        -- Test 4: �H���t�׼Ҧ�
        report "Test 4: Random speed";
        i_speed_switch <= '1';
        i_right_button <= '1';
        wait for 100 ns;
        i_right_button <= '0';
        wait for 2000 ns;
        
        report "Tests done";
        test_done <= true;
        wait;
    end process;

end Behavioral;